module test;
  initial begin
    $display("Hello, Icarus!");
    $finish;
  end
endmodule